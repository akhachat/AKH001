module PEM00X(
);
endmodule
